


G1  1 2 4 3 VCCS_K
R1  4 3 R
v1  1 2 5

.end
