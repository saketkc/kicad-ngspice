


G1  3 4 1 2 VCCS_K
R1  4 3 R
v1  1 2 5


.end
