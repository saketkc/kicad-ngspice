* EESchema Netlist Version 1.1 (Spice format) creation date: Thursday 29 September 2011 08:12:07 PM IST


K1_L1_L2  0.87
R2  0 3 100
R1  2 1 100
L2  0 3 1m
L1  2 0 1m

.end
