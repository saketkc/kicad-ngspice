* EESchema Netlist Version 1.1 (Spice format) creation date: Tuesday 04 October 2011 07:17:27 PM IST


v2  2 0 sin(0 5 1khz)
R1  4 0 200
v1  1 0 15
m1  1 2 4 1 MOSFET_P 
m2  4 2 0 0 MOSFET_N 

.end

