* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 21 November 2011 02:11:51 AM IST

.MODEL TR NPN(BF=140 CJC=20pf CJE=20pf IS=1E-16 VJE =0.7)

v4  7 1 0
R4  7 0 3.9k
Q1  6 1 2 TR
R3  2 0 1.5k
v3  4 5 0
v1  4 0 22
R1  4 7 39k
R2  5 6 10k

.tran 1ms 100ms

.control
run
.endc

.end
