* EESchema Netlist Version 1.1 (Spice format) creation date: Thursday 29 September 2011 08:55:39 PM IST


R1  1 4 R
v  3 2 5
E1  3 2 1 4 VCVS_K1

.end
