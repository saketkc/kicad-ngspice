* EESchema Netlist Version 1.1 (Spice format) creation date: Saturday 01 October 2011 12:59:44 PM IST


v1  3 0 AC
R1  2 0 1k
C1  2 3 3.3nf

.end
