* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 03 October 2011 04:01:36 PM IST


F1  6 1 vc 5
vc1  2 3 0
R3  6 0 47
R1  5 3 100
R2  1 0 32
v1  2 0 10

.end
